library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.std_logic_arith.ALL;

--                       General timing
--          Screen refresh rate |   60 Hz
--          Vertical refresh    |   31.46875 kHz
--          Pixel freq          |   25.175 MHz

--                  Horizontal timing (line)
--          Scanline part |	Pixels | Time [µs]
--          Visible area  |  640   |  25.422045680238
--          Front porch	  |   16   |  0.63555114200596
--          Sync pulse	  |   96   |  3.8133068520357
--          Back porch	  |   48   |  1.9066534260179
--          Whole line	  |  800   |  31.777557100298

--                  Vertical timing (frame)
--          Scanline part |	Pixels | Time [µs]
--          Visible area  |  480   |  15.253227408143
--          Front porch	  |   10   |  0.31777557100298
--          Sync pulse	  |   2    |  0.063555114200596
--          Back porch	  |   33   |  1.0486593843098
--          Whole line	  |  525   |  16.683217477656

entity VGA_Sync is
    --  Generic ( );
    --  Port ( );
    port(
        -- Inputs
        clk   : in std_logic;
        -- Outputs
        rgb   : out std_logic_vector(11 downto 0);
        HSync : out std_logic;
        VSync : out std_logic
        
    );
end VGA_Sync;

-- Bit    7  6  5  4  3  2  1  0
-- Data   R  R  R  G  G  G  B  B

architecture rtl of VGA_Sync is

    -- Declarative zone of VHDL

    --Horizontal Synchronization Constants
    constant Active_Cols: integer:= 640;
    constant Front_HPorch: integer:= 16;
    constant SP_H: integer:= 96;
    constant Back_HPorch: integer:= 48;
    constant Total_Cols: integer:= Active_Cols + Front_HPorch + SP_H + Back_HPorch; --800 in total
    
    --Vertical Synchronization Constants
    constant Active_Rows: integer:= 480;
    constant Front_VPorch: integer:= 10;
    constant SP_V: integer:= 2;
    constant Back_Vporch: integer:= 33;
    constant Total_Rows: integer:= Active_Rows + Front_VPorch + SP_V + Back_Vporch; --525 in total
    
    signal vPos : integer range 0 to Total_Rows - 1 := 0; -- They go to all display 800 x 525
    signal hPos : integer range 0 to Total_Cols - 1 := 0;
    
    signal videoOn : std_logic := '0';
    
    --Defitions of the bitmaps for different images, they will be stored in the ROM 

    type BITMAP is array (0 to 164) of std_logic_vector(0 to 199);
    signal logo: BITMAP := 
            ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111111111111111111111111",
             "11111111111111111111111111111111111000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111111",
             "11111111111111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000000000000000000000000000000001111111111111111111111111111111",
             "11111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111",
             "11111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111",
             "11111111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000011111111111111111111111111",
             "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
             "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
             "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
             "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
             "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
             "11111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111",
             "11111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111",
             "11111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111",
             "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111",
             "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111",
             "11111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111",
             "11111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111",
             "11111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111",
             "11111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
             "11111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
             "11111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
             "11111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
             "11111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
             "11111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
             "11111111111000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
             "11111111111000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
             "11111111111000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
             "11111111111110000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
             "11111111111110000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
             "11111111111111000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
             "11111111111111000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
             "11111111111111100000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
             "11111111111111100000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111",
             "11111111111111110000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111",
             "11111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111",
             "11111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111",
             "11111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111",
             "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111",
             "11111111111111111110000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111",
             "11111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111",
             "11111111111111111111000000000000000000000000000000000000000000000000000000000000000000011111001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111",
             "11111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111100011111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111",
             "11111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111100000111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111",
             "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000000111100000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
             "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000000011110000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
             "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011110000000001111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
             "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011110000000000011111111000000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
             "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111000000000001111111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
             "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111000000000000011111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
             "11111111111111111111111111100000000000000000000000000000000000000000000000000000000001111111111000000000000000111111110000000000000000000000000000000000000000000000000000000001111111111111111111111111",
             "11111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111111111111",
             "11111111111111111111111111111000000000000000000000000000000000000000000000000000001111111100111000000000000000000111111111000000000000000000000000000000000000000000000000000011111111111111111111111111",
             "11111111111111111111111111111100000000000000000000000000000000000000000000000000111111110001111000000000000000000001111111100000000000000000000000000000000000000000000000000111111111111111111111111111",
             "11111111111111111111111111111110000000000000000000000000000000000000000000000011111111000001111000000000000000000000111111111000000000000000000000000000000000000000000000001111111111111111111111111111",
             "11111111111111111111111111111111000000000000000000000000000000000000000000000111111110000001111000000000000000000000001111111110000000000000000000000000000000000000000000011111111111111111111111111111",
             "11111111111111111111111111111111100000000000000000000000000000000000000000011111111000000001111000000000000000000000000011111111000000000000000000000000000000000000000000111111111111111111111111111111",
             "11111111111111111111111111111111110000000000000000000000000000000000000001111111100000000001110000000000000000000000000001111111110000000000000000000000000000000000000001111111111111111111111111111111",
             "11111111111111111111111111111111111000000000000000000000000000000000000011111110000000000011110000000000000000000000000000011111111100000000000000000000000000000000000111111111111111111111111111111111",
             "11111111111111111111111111111111111100000000000000000000000000000000001111111100000000000011110000000000000000000000000000000111111110000000000000000000000000000000001111111111111111111111111111111111",
             "11111111111111111111111111111111111111000000000000000000000000000000111111110000000000000111110000000000000000000000000000000001111111100000000000000000000000000000011111111111111111111111111111111111",
             "11111111111111111111111111111111111111100000000000000000000000000011111111000000000000000111100000000000000000000000000000000000111111111000000000000000000000000001111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111000000000000000000000000111111110000000000000001111100000000000000000000000000000000000001111111100000000000000000000000111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111110000000000000000000011111111000000000000000001111000000000000000000000000000000000000000011111111000000000000000000011111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111000000000000000001111111100000000000000000011111000000000000000000000000000000000000000001111111110000000000000001111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111000000000000111111111000000000000000000011110000000000000000000000000000000000000000000011111111110000000001111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111000000111111111111111111000000000000111110000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111110000001111100000000000000000000000111110000001111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111100000011111100000000000000000000001111111000001111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111000000111111100000000000000000000001111111000000111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111000001111111110000000000000000000001111111100000011111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111110000001111111100000000000000000000001111111110000011111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000000000000000000000111111111000001111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111000000111111111000000000000000000000000111111111000000111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111000001111111111000000000000000000000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111110000001111111110000000000001100000000000001111111110000011111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000000000001110000000000001111111110000001111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111000000111111111100000000000011110000000000000111111111000000111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111000000111111111000000000000111111000000000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111110000001111111110000000000000111111100000000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111100000011111111100000000000001111111100000000000001111111110000001111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111100000011111111100000000000001111111110000000000000111111111000000111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111000000111111111000000000000011111111111000000000000111111111100000111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111110000001111111110000000000000111111111111000000000000011111111100000011111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111100000001111111110000000000000111111111111100000000000001111111110000001111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111100000001111111100000000000001111111111111110000000000000111111110000000111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111000000001111111000000000000011111111111111110000000000000111111110000000111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111110000000000111110000000000000011111111111111111000000000000011111100000000011111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111110000000000011100000000000000111111111111111111100000000000000110000000000001111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000011111111111111111111110000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

    type BITMAP1 is array (0 to 60) of std_logic_vector(0 to 299);
    signal message : BITMAP1 :=
               ("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011001111111111111",
                "111100000000011111111100000000011111111111111000000000111111111111111000000000111111111000000000111111111111111111111111111111100000000011111100000000011111100000000011111111111111100000000011111111111111111111111000000000001111111111111111111111111111111111111111111111111111111011001100111111111111",
                "111101101010001111111101001010001111111111100011111110001111111111111001010110011111111011010100011111111111111111111111111111101101010001111101101011001111101001010001111111111110001111111000111111111111111111110011111111100011111111111111111111111111111111111111111111111111111000110110111111111111",
                "111101101010000111111101001010000111111110011110000011100111111111111001010110001111111011010100001111111111111111111111111111101101010000111101101011000111101001010000111111111001110000001110011111111111111111001110000000011001111111111111111111111111111111111111111111111111111010011010011111111111",
                "111101101010000011111101001010000011111100110001111100011001111111111001010110000111111011010100000111111111111111111111111111101101010000011101101011000011101001010000011111110011000111110001100111111111111110011001111111000100111111111111111111111111111111111111111111111111111001001001001111111111",
                "111101101010000001111101001010000011111001100111000111001100111111111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011111100110011100011100110011111111111100110111000001110010011111111111111111111111111111111111111111111111111000100101000111111111",
                "111101101010000001111101001010000011111011011000000000110110111111111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011111101101100000000011011011111111111101101100011100011001001111111111111111111111111111111111111111111111111100110100100011111111",
                "111101101010000001111101001010000011110110110011111110011011011111111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011111011011001111111001101101111111111011011001110111100100100111111111111111111111111111111111111111111111111110010100100001111111",
                "111101101010000001111101001010000011100100100100000001001001001111111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011110010010010000000100100100111111111010010010000000110110110011111111111111111111111111111111111111111111111111010010100001111111",
                "111101101010000001111101001010000011101101001000000000100101100111111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011110110100100000000010010110011111110010100100000000011010010001111111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011101001010000000000010100100011111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011110100101000000000001010010001111110100101000000000001001010000111111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011101010010000000000010010100001111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011110101001000000000001001010000111110100101000000000001001010000111111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011001010010000000000011010100000111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101001000000000001101010000111110101001000000000000101011000011111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011001010010000000111011010100000111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101001000000011101101010000011110101001000000011100101011000011111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011001010010000001111011010110000111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000000111101101010000011110101001000000111100101011000011111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011001010010000011111011010110000111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000011110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111100101011000001111101001010000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111100101001000001111101010010000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111110101101000001111001010010000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111110100100100001110010010100000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111110010110011000000100100100000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111111011011001111111001001000000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111110001111111111111010010100000111111",
                "111111001001110000000010011000000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111000100011111111111010010100000111111",
                "111111100100011110111100110000000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111011111011111111111010010100000111111",
                "111111110011000111100001100000000111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111110010001001111111111010010100000111111",
                "111111111001110001000110000000000111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111110110101000111111111010010100000111111",
                "111111111100001101011000000000001111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111110010001000011111111010010100000111111",
                "111111111110001101010000000000001111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111011111000001111111010010100000111111",
                "111111111111001101010000000000011111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111000100000000111111010010100000111111",
                "111111111111101101010000000000111111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111100000000000111111010010100000111111",
                "111111111111101101010000000011111111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111000000000111111010010100000111111",
                "111111111111101101010000001111111111001010010000011111011010100000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111100000001111111010010100000111111",
                "111111111111101101010000001111111111001010010000011111011010100000011001010010000011111010010100000011111111111111111111111111101101010000001101101011000001101001010000011100101001000001111101101010000001110101001000001111100101011000001111111111111111111111111111111110000001111111010010100000111111",
                "111111111111101101010000001111111111101010010000011111010010100000011001010010000011111010010100000011111111111111111111111111101101010000001101001001000001101001010000011110101001000001111101001010000001110101001000001111100101011000001111111111111111111111111111111111000111111111010010100000111111",
                "111111111111101101010000001111111111101001010000011111010110100000011101011010000011110010100100000011111111111111111111111111100101001000001001011101000001101001010000011110100101000001111101011010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111111111111101101010000001111111111101101001000011110010100100000011101101001000011100100100100000011111111111111111111111111100101001000000011011101100001001011010000011110110100100001111001010010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111111111111101101010000001111111111100100101100010000101101100000011100101101100000001101101000000011111111111111111111111111110100100100000110110110100000010010010000011110010010110001000010110100000001110101001000001111100101011000001111111111111111111111111111110001111111111111010010100000111111",
                "111111111111101101010000001111111111110110110111000011001001000000011110110110011111111001001000000111111111111111111111111111110100110011111100100010011111100110100000011111011010011100001100100100000001110101001000001111100101011000001111111111111111111111111111000100011111111111010110100000111111",
                "111111111111101101010000001111111111110010011001111100110010000000111110010011000111000110010000000111111111111111111111111111110010011000110001100011000110001100100000011111001001100111110011001000000011110101001000001111100101011000001111111111111111111111111111011111011111111110010100100000111111",
                "111111111111101101010000001111111111111001001100000001100110000000111111001001110000011100100000000111111111111111111111111111111011001110000110011101110000111001000000011111100100110000000110011000000011110101001000001111100101011000001111111111111111111111111110010001001111111100100101000000111111",
                "111111111111101101010000001111111111111100100011111111001100000000111111100110011111110001000000000111111111111111111111111111111101100011111100110100011111100010000000011111110010001111111100110000000011110101001000001111100101011000001111111111111111111111111110110101000111111001001001000000111111",
                "111111111111101101010000001111111111111110011000000000110000000000111111110011000000000110000000001111111111111111111111111111111100111000000001100011000000001100000000011111111001100000000011000000000111110101001000001111100101011000001111111111111111111111111110010001000011111010011011000000111111",
                "111111111111101101010000001111111111111111001111000111100000000001111111111000111111111000000000001111111111111111111111111111111111001111111110000000111111111000000000111111111100111100011110000000000111110101001000001111100101011000001111111111111111111111111111011110000001111000110110000000111111",
                "111111111111100001000000001111111111111111100001111100000000000011111111111100000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000111111111110000111110000000000001111110100000000001111100001000000001111111111111111111111111111000000000000111011101100000000111111",
                "111111111111100000000000001111111111111111110000000000000000000011111111111110000000000000000000111111111111111111111111111111111111110000000000000000000000000000000001111111111111000000000000000000011111110000000000001111110000000000001111111111111111111111111111110000000000111010011000000001111111",
                "111111111111110000000000001111111111111111111000000000000000000111111111111111000000000000000001111111111111111111111111111111111111111000000000000000000000000000000011111111111111100000000000000000011111111000000000001111111000000000001111111111111111111111111111111000000000111001110000000001111111",
                "111111111111111000000000001111111111111111111100000000000000011111111111111111100000000000000011111111111111111111111111111111111111111100000000000000110000000000000111111111111111110000000000000001111111111100000000001111111100000000001111111111111111111111111111111100000001111011000000000011111111",
                "111111111111111100000000001111111111111111111111000000000000111111111111111111111000000000001111111111111111111111111111111111111111111110000000000011111000000000001111111111111111111100000000000011111111111110000000001111111110000000001111111111111111111111111111111110000001111000000000000011111111",
                "111111111111111111000000011111111111111111111111110000000111111111111111111111111111000001111111111111111111111111111111111111111111111111110000011111111111000001111111111111111111111111000000011111111111111111000000001111111111000000001111111111111111111111111111111111000111111000000000000111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000001111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
            
    signal logoVisible : boolean := false;   
    signal logoColor : std_logic_vector(11 downto 0) := "000010101110";
    
    signal messageVisible : boolean := false;
    signal messageColor : std_logic_vector(11 downto 0) := "001110100010";
    
begin
       
   -- Out signal assigment
   HSync <= '1' when hPos < Active_Cols + Front_HPorch or hPos > Active_Cols + Front_HPorch + SP_H  else '0'; -- Add Front and Back porch for image to be centered
   VSync <= '1' when vPos < Active_Rows + Front_VPorch or vPos > Active_Rows + Front_VPorch + SP_V  else '0'; -- Add Front and Back porch for image to be centered

   videoOn <= '1' when hPos < Active_Cols and vPos < Active_Rows else '0'; -- Active Area
   
   logoVisible <= (vPos >= (Active_Rows / 2) -  45) and (vPos < (Active_Rows / 2) + 120) and
                  (hPos >= (Active_Cols / 2) - 100) and (hPos < (Active_Cols / 2) + 100) and
                  logo(vPos - ((Active_Rows / 2) - 45))(hPos - ((Active_Cols / 2) - 100)) = '0';
                  
   messageVisible <= (vPos >= (Active_Rows / 4) -  30) and (vPos < (Active_Rows / 4) +  31) and
                     (hPos >= (Active_Cols / 2) - 150) and (hPos < (Active_Cols / 2) + 150) and
                     message(vPos - ((Active_Rows / 4) -  30))(hPos - ((Active_Cols / 2) - 150)) = '0';
   
   rgb(11 downto 0) <= logoColor(11 downto 0)    when logoVisible = true    and videoOn = '1' else
                       messageColor(11 downto 0) when messageVisible = true and videoOn = '1' else
                       (others => '0');
    
   Sync_proc : process(clk) is
   begin
    if rising_edge(clk) then
        if hPos = Total_Cols - 1 then
            if vPos = Total_Rows - 1 then
                vPos <= 0;
            else
                vPos <= vPos + 1;
            end if;
            hPos <= 0;
        else
            hPos <= hPos + 1;
        end if;
    end if;
   end process Sync_proc;

end rtl;
